`default_nettype none
module ksatask2(CLOCK_50, KEY, SW, LEDR, HEX5, HEX4, HEX3, HEX2, HEX1, HEX0);

input CLOCK_50;
input [3:0] KEY;
input [9:0] SW;
output [9:0] LEDR;
output [6:0] HEX5, HEX4, HEX3, HEX2, HEX1, HEX0;

//hex display inputs
reg [3:0]inHEX0;
reg [3:0]inHEX1;
reg [3:0]inHEX2;
reg [3:0]inHEX3;
reg [3:0]inHEX4;
reg [3:0]inHEX5;
//reset
assign reset = ~KEY[3];
assign CLK_50M = CLOCK_50;

//Seven Segment 
SevenSegmentDisplayDecoder U0(HEX0, inHEX0);
SevenSegmentDisplayDecoder U1(HEX1, inHEX1);
SevenSegmentDisplayDecoder U2(HEX2, inHEX2);
SevenSegmentDisplayDecoder U3(HEX3, inHEX3);
SevenSegmentDisplayDecoder U4(HEX4, inHEX4);
SevenSegmentDisplayDecoder U5(HEX5, inHEX5);
wire [7:0] address;
wire [7:0] i ;
wire [7:0] data;
wire [7:0]q;
wire wren;

s_memory s1 (
	.address(address),
	.clock(CLOCK_50),
	.data(data),
	.wren(wren),
	.q(q));

reg [3:0] state;

reg [3:0] initial_state = 4'b0;

	always_ff @(posedge CLK_50M, posedge reset) 
	if (reset) begin
		state <= initial_state;
		i <= 8'b0;
	end 
	else begin
		case (state)
			initial_state: begin
				LEDR[9:0] = 10'b0;
				state <= s_init_task1;
			end 
			
			s_init_task1: begin 
				i <= 8'b0;
				state <= s_increment;
				wren <= 1'b1;
			end 
			
			s_increment: begin
				address <= i[7:0];
				data <= i[7:0];
				wren <= 1'b1;
				i <= i + 8'd1;
				if (i == 255) begin
					state <= s_init_task2a;
				end
				else state <= s_increment;
endmodule

